architecture ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sig3 is

end entity;

architecture rtl of sig3 is
end architecture;
