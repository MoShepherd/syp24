library ieee;
use ieee.std_logic_1164.all;

package mem_buffer is
  constant address_size : integer := 10;  -- ram_adddress breite
  type mem_type is array (0 to (2**address_size)-1) of std_logic_vector(15 downto 0);

  constant mem_buffer_image : mem_type := (
      0  => "1010101010101010",
      1  => "1010101010101010",
      2  => "1010101010101010",
      3  => "1010101010101010",
      4  => "1010101010101010",
      5  => "1010101010101010",
      6  => "1010101010101010",
      7  => "1010101010101010",
      8  => "1010101010101010",
      9  => "1010101010101010",
     10  => "1010101010101010",
     11  => "1010101010101010",
     12  => "1010101010101010",
     13  => "1010101010101010",
     14  => "1010101010101010",
     15  => "1010101010101010",
     16  => "1010101010101010",
     17  => "1010101010101010",
     18  => "1010101010101010",
     19  => "1010101010101010",
     20  => "1010101010101010",
     21  => "1010101010101010",
     22  => "1010101010101010",
     23  => "1010101010101010",
     24  => "1010101010101010",
     25  => "1010101010101010",
     26  => "1010101010101010",
     27  => "1010101010101010",
     28  => "1010101010101010",
     29  => "1010101010101010",
     30  => "1010101010101010",
     31  => "1010101010101010",
     32  => "1010101010101010",
     33  => "1010101010101010",
     34  => "1010101010101010",
     35  => "1010101010101010",
     36  => "1010101010101010",
     37  => "1010101010101010",
     38  => "1010101010101010",
     39  => "1010101010101010",
     40  => "1010101010101010",
     41  => "1010101010101010",
     42  => "1010101010101010",
     43  => "1010101010101010",
     44  => "1010101010101010",
     45  => "1010101010101010",
     46  => "1010101010101010",
     47  => "1010101010101010",
     48  => "1010101010101010",
     49  => "1010101010101010",
     50  => "1010101010101010",
     51  => "1010101010101010",
     52  => "1010101010101010",
     53  => "1010101010101010",
     54  => "1010101010101010",
     55  => "1010101010101010",
     56  => "1010101010101010",
     57  => "1010101010101010",
     58  => "1010101010101010",
     59  => "1010101010101010",
     60  => "1010101010101010",
     61  => "1010101010101010",
     62  => "1010101010101010",
     63  => "1010101010101010",
     64  => "1010101010101010",
     65  => "1010101010101010",
     66  => "1010101010101010",
     67  => "1010101010101010",
     68  => "1010101010101010",
     69  => "1010101010101010",
     70  => "1010101010101010",
     71  => "1010101010101010",
     72  => "1010101010101010",
     73  => "1010101010101010",
     74  => "1010101010101010",
     75  => "1010101010101010",
     76  => "1010101010101010",
     77  => "1010101010101010",
     78  => "1010101010101010",
     79  => "1010101010101010",
     80  => "1010101010101010",
     81  => "1010101010101010",
     82  => "1010101010101010",
     83  => "1010101010101010",
     84  => "1010101010101010",
     85  => "1010101010101010",
     86  => "1010101010101010",
     87  => "1010101010101010",
     88  => "1010101010101010",
     89  => "1010101010101010",
     90  => "1010101010101010",
     91  => "1010101010101010",
     92  => "1010101010101010",
     93  => "1010101010101010",
     94  => "1010101010101010",
     95  => "1010101010101010",
     96  => "1010101010101010",
     97  => "1010101010101010",
     98  => "1010101010101010",
     99  => "1010101010101010",
    100  => "1010101010101010",
    101  => "1010101010101010",
    102  => "1010101010101010",
    103  => "1010101010101010",
    104  => "1010101010101010",
    105  => "1010101010101010",
    106  => "1010101010101010",
    107  => "1010101010101010",
    108  => "1010101010101010",
    109  => "1010101010101010",
    110  => "1010101010101010",
    111  => "1010101010101010",
    112  => "1010101010101010",
    113  => "1010101010101010",
    114  => "1010101010101010",
    115  => "1010101010101010",
    116  => "1010101010101010",
    117  => "1010101010101010",
    118  => "1010101010101010",
    119  => "1010101010101010",
    120  => "1010101010101010",
    121  => "1010101010101010",
    122  => "1010101010101010",
    123  => "1010101010101010",
    124  => "1010101010101010",
    125  => "1010101010101010",
    126  => "1010101010101010",
    127  => "1010101010101010",
    128  => "1010101010101010",
    129  => "1010101010101010",
    130  => "1010101010101010",
    131  => "1010101010101010",
    132  => "1010101010101010",
    133  => "1010101010101010",
    134  => "1010101010101010",
    135  => "1010101010101010",
    136  => "1010101010101010",
    137  => "1010101010101010",
    138  => "1010101010101010",
    139  => "1010101010101010",
    140  => "1010101010101010",
    141  => "1010101010101010",
    142  => "1010101010101010",
    143  => "1010101010101010",
    144  => "1010101010101010",
    145  => "1010101010101010",
    146  => "1010101010101010",
    147  => "1010101010101010",
    148  => "1010101010101010",
    149  => "1010101010101010",
    150  => "1010101010101010",
    151  => "1010101010101010",
    152  => "1010101010101010",
    153  => "1010101010101010",
    154  => "1010101010101010",
    155  => "1010101010101010",
    156  => "1010101010101010",
    157  => "1010101010101010",
    158  => "1010101010101010",
    159  => "1010101010101010",
    160  => "1010101010101010",
    161  => "1010101010101010",
    162  => "1010101010101010",
    163  => "1010101010101010",
    164  => "1010101010101010",
    165  => "1010101010101010",
    166  => "1010101010101010",
    167  => "1010101010101010",
    168  => "1010101010101010",
    169  => "1010101010101010",
    170  => "1010101010101010",
    171  => "1010101010101010",
    172  => "1010101010101010",
    173  => "1010101010101010",
    174  => "1010101010101010",
    175  => "1010101010101010",
    176  => "1010101010101010",
    177  => "1010101010101010",
    178  => "1010101010101010",
    179  => "1010101010101010",
    180  => "1010101010101010",
    181  => "1010101010101010",
    182  => "1010101010101010",
    183  => "1010101010101010",
    184  => "1010101010101010",
    185  => "1010101010101010",
    186  => "1010101010101010",
    187  => "1010101010101010",
    188  => "1010101010101010",
    189  => "1010101010101010",
    190  => "1010101010101010",
    191  => "1010101010101010",
    192  => "1010101010101010",
    193  => "1010101010101010",
    194  => "1010101010101010",
    195  => "1010101010101010",
    196  => "1010101010101010",
    197  => "1010101010101010",
    198  => "1010101010101010",
    199  => "1010101010101010",
    200  => "1010101010101010",
    201  => "1010101010101010",
    202  => "1010101010101010",
    203  => "1010101010101010",
    204  => "1010101010101010",
    205  => "1010101010101010",
    206  => "1010101010101010",
    207  => "1010101010101010",
    208  => "1010101010101010",
    209  => "1010101010101010",
    210  => "1010101010101010",
    211  => "1010101010101010",
    212  => "1010101010101010",
    213  => "1010101010101010",
    214  => "1010101010101010",
    215  => "1010101010101010",
    216  => "1010101010101010",
    217  => "1010101010101010",
    218  => "1010101010101010",
    219  => "1010101010101010",
    220  => "1010101010101010",
    221  => "1010101010101010",
    222  => "1010101010101010",
    223  => "1010101010101010",
    224  => "1010101010101010",
    225  => "1010101010101010",
    226  => "1010101010101010",
    227  => "1010101010101010",
    228  => "1010101010101010",
    229  => "1010101010101010",
    230  => "1010101010101010",
    231  => "1010101010101010",
    232  => "1010101010101010",
    233  => "1010101010101010",
    234  => "1010101010101010",
    235  => "1010101010101010",
    236  => "1010101010101010",
    237  => "1010101010101010",
    238  => "1010101010101010",
    239  => "1010101010101010",
    240  => "1010101010101010",
    241  => "1010101010101010",
    242  => "1010101010101010",
    243  => "1010101010101010",
    244  => "1010101010101010",
    245  => "1010101010101010",
    246  => "1010101010101010",
    247  => "1010101010101010",
    248  => "1010101010101010",
    249  => "1010101010101010",
    250  => "1010101010101010",
    251  => "1010101010101010",
    252  => "1010101010101010",
    253  => "1010101010101010",
    254  => "1010101010101010",
    255  => "1010101010101010",
    256  => "1010101010101010",
    257  => "1010101010101010",
    258  => "1010101010101010",
    259  => "1010101010101010",
    260  => "1010101010101010",
    261  => "1010101010101010",
    262  => "1010101010101010",
    263  => "1010101010101010",
    264  => "1010101010101010",
    265  => "1010101010101010",
    266  => "1010101010101010",
    267  => "1010101010101010",
    268  => "1010101010101010",
    269  => "1010101010101010",
    270  => "1010101010101010",
    271  => "1010101010101010",
    272  => "1010101010101010",
    273  => "1010101010101010",
    274  => "1010101010101010",
    275  => "1010101010101010",
    276  => "1010101010101010",
    277  => "1010101010101010",
    278  => "1010101010101010",
    279  => "1010101010101010",
    280  => "1010101010101010",
    281  => "1010101010101010",
    282  => "1010101010101010",
    283  => "1010101010101010",
    284  => "1010101010101010",
    285  => "1010101010101010",
    286  => "1010101010101010",
    287  => "1010101010101010",
    288  => "1010101010101010",
    289  => "1010101010101010",
    290  => "1010101010101010",
    291  => "1010101010101010",
    292  => "1010101010101010",
    293  => "1010101010101010",
    294  => "1010101010101010",
    295  => "1010101010101010",
    296  => "1010101010101010",
    297  => "1010101010101010",
    298  => "1010101010101010",
    299  => "1010101010101010",
    300  => "1010101010101010",
    301  => "1010101010101010",
    302  => "1010101010101010",
    303  => "1010101010101010",
    304  => "1010101010101010",
    305  => "1010101010101010",
    306  => "1010101010101010",
    307  => "1010101010101010",
    308  => "1010101010101010",
    309  => "1010101010101010",
    310  => "1010101010101010",
    311  => "1010101010101010",
    312  => "1010101010101010",
    313  => "1010101010101010",
    314  => "1010101010101010",
    315  => "1010101010101010",
    316  => "1010101010101010",
    317  => "1010101010101010",
    318  => "1010101010101010",
    319  => "1010101010101010",
    320  => "1010101010101010",
    321  => "1010101010101010",
    322  => "1010101010101010",
    323  => "1010101010101010",
    324  => "1010101010101010",
    325  => "1010101010101010",
    326  => "1010101010101010",
    327  => "1010101010101010",
    328  => "1010101010101010",
    329  => "1010101010101010",
    330  => "1010101010101010",
    331  => "1010101010101010",
    332  => "1010101010101010",
    333  => "1010101010101010",
    334  => "1010101010101010",
    335  => "1010101010101010",
    336  => "1010101010101010",
    337  => "1010101010101010",
    338  => "1010101010101010",
    339  => "1010101010101010",
    340  => "1010101010101010",
    341  => "1010101010101010",
    342  => "1010101010101010",
    343  => "1010101010101010",
    344  => "1010101010101010",
    345  => "1010101010101010",
    346  => "1010101010101010",
    347  => "1010101010101010",
    348  => "1010101010101010",
    349  => "1010101010101010",
    350  => "1010101010101010",
    351  => "1010101010101010",
    352  => "1010101010101010",
    353  => "1010101010101010",
    354  => "1010101010101010",
    355  => "1010101010101010",
    356  => "1010101010101010",
    357  => "1010101010101010",
    358  => "1010101010101010",
    359  => "1010101010101010",
    360  => "1010101010101010",
    361  => "1010101010101010",
    362  => "1010101010101010",
    363  => "1010101010101010",
    364  => "1010101010101010",
    365  => "1010101010101010",
    366  => "1010101010101010",
    367  => "1010101010101010",
    368  => "1010101010101010",
    369  => "1010101010101010",
    370  => "1010101010101010",
    371  => "1010101010101010",
    372  => "1010101010101010",
    373  => "1010101010101010",
    374  => "1010101010101010",
    375  => "1010101010101010",
    376  => "1010101010101010",
    377  => "1010101010101010",
    378  => "1010101010101010",
    379  => "1010101010101010",
    380  => "1010101010101010",
    381  => "1010101010101010",
    382  => "1010101010101010",
    383  => "1010101010101010",
    384  => "1010101010101010",
    385  => "1010101010101010",
    386  => "1010101010101010",
    387  => "1010101010101010",
    388  => "1010101010101010",
    389  => "1010101010101010",
    390  => "1010101010101010",
    391  => "1010101010101010",
    392  => "1010101010101010",
    393  => "1010101010101010",
    394  => "1010101010101010",
    395  => "1010101010101010",
    396  => "1010101010101010",
    397  => "1010101010101010",
    398  => "1010101010101010",
    399  => "1010101010101010",
    400  => "1010101010101010",
    401  => "1010101010101010",
    402  => "1010101010101010",
    403  => "1010101010101010",
    404  => "1010101010101010",
    405  => "1010101010101010",
    406  => "1010101010101010",
    407  => "1010101010101010",
    408  => "1010101010101010",
    409  => "1010101010101010",
    410  => "1010101010101010",
    411  => "1010101010101010",
    412  => "1010101010101010",
    413  => "1010101010101010",
    414  => "1010101010101010",
    415  => "1010101010101010",
    416  => "1010101010101010",
    417  => "1010101010101010",
    418  => "1010101010101010",
    419  => "1010101010101010",
    420  => "1010101010101010",
    421  => "1010101010101010",
    422  => "1010101010101010",
    423  => "1010101010101010",
    424  => "1010101010101010",
    425  => "1010101010101010",
    426  => "1010101010101010",
    427  => "1010101010101010",
    428  => "1010101010101010",
    429  => "1010101010101010",
    430  => "1010101010101010",
    431  => "1010101010101010",
    432  => "1010101010101010",
    433  => "1010101010101010",
    434  => "1010101010101010",
    435  => "1010101010101010",
    436  => "1010101010101010",
    437  => "1010101010101010",
    438  => "1010101010101010",
    439  => "1010101010101010",
    440  => "1010101010101010",
    441  => "1010101010101010",
    442  => "1010101010101010",
    443  => "1010101010101010",
    444  => "1010101010101010",
    445  => "1010101010101010",
    446  => "1010101010101010",
    447  => "1010101010101010",
    448  => "1010101010101010",
    449  => "1010101010101010",
    450  => "1010101010101010",
    451  => "1010101010101010",
    452  => "1010101010101010",
    453  => "1010101010101010",
    454  => "1010101010101010",
    455  => "1010101010101010",
    456  => "1010101010101010",
    457  => "1010101010101010",
    458  => "1010101010101010",
    459  => "1010101010101010",
    460  => "1010101010101010",
    461  => "1010101010101010",
    462  => "1010101010101010",
    463  => "1010101010101010",
    464  => "1010101010101010",
    465  => "1010101010101010",
    466  => "1010101010101010",
    467  => "1010101010101010",
    468  => "1010101010101010",
    469  => "1010101010101010",
    470  => "1010101010101010",
    471  => "1010101010101010",
    472  => "1010101010101010",
    473  => "1010101010101010",
    474  => "1010101010101010",
    475  => "1010101010101010",
    476  => "1010101010101010",
    477  => "1010101010101010",
    478  => "1010101010101010",
    479  => "1010101010101010",
    480  => "1010101010101010",
    481  => "1010101010101010",
    482  => "1010101010101010",
    483  => "1010101010101010",
    484  => "1010101010101010",
    485  => "1010101010101010",
    486  => "1010101010101010",
    487  => "1010101010101010",
    488  => "1010101010101010",
    489  => "1010101010101010",
    490  => "1010101010101010",
    491  => "1010101010101010",
    492  => "1010101010101010",
    493  => "1010101010101010",
    494  => "1010101010101010",
    495  => "1010101010101010",
    496  => "1010101010101010",
    497  => "1010101010101010",
    498  => "1010101010101010",
    499  => "1010101010101010",
    500  => "1010101010101010",
    501  => "1010101010101010",
    502  => "1010101010101010",
    503  => "1010101010101010",
    504  => "1010101010101010",
    505  => "1010101010101010",
    506  => "1010101010101010",
    507  => "1010101010101010",
    508  => "1010101010101010",
    509  => "1010101010101010",
    510  => "1010101010101010",
    511  => "1010101010101010",
    512  => "1010101010101010",
    513  => "1010101010101010",
    514  => "1010101010101010",
    515  => "1010101010101010",
    516  => "1010101010101010",
    517  => "1010101010101010",
    518  => "1010101010101010",
    519  => "1010101010101010",
    520  => "1010101010101010",
    521  => "1010101010101010",
    522  => "1010101010101010",
    523  => "1010101010101010",
    524  => "1010101010101010",
    525  => "1010101010101010",
    526  => "1010101010101010",
    527  => "1010101010101010",
    528  => "1010101010101010",
    529  => "1010101010101010",
    530  => "1010101010101010",
    531  => "1010101010101010",
    532  => "1010101010101010",
    533  => "1010101010101010",
    534  => "1010101010101010",
    535  => "1010101010101010",
    536  => "1010101010101010",
    537  => "1010101010101010",
    538  => "1010101010101010",
    539  => "1010101010101010",
    540  => "1010101010101010",
    541  => "1010101010101010",
    542  => "1010101010101010",
    543  => "1010101010101010",
    544  => "1010101010101010",
    545  => "1010101010101010",
    546  => "1010101010101010",
    547  => "1010101010101010",
    548  => "1010101010101010",
    549  => "1010101010101010",
    550  => "1010101010101010",
    551  => "1010101010101010",
    552  => "1010101010101010",
    553  => "1010101010101010",
    554  => "1010101010101010",
    555  => "1010101010101010",
    556  => "1010101010101010",
    557  => "1010101010101010",
    558  => "1010101010101010",
    559  => "1010101010101010",
    560  => "1010101010101010",
    561  => "1010101010101010",
    562  => "1010101010101010",
    563  => "1010101010101010",
    564  => "1010101010101010",
    565  => "1010101010101010",
    566  => "1010101010101010",
    567  => "1010101010101010",
    568  => "1010101010101010",
    569  => "1010101010101010",
    570  => "1010101010101010",
    571  => "1010101010101010",
    572  => "1010101010101010",
    573  => "1010101010101010",
    574  => "1010101010101010",
    575  => "1010101010101010",
    576  => "1010101010101010",
    577  => "1010101010101010",
    578  => "1010101010101010",
    579  => "1010101010101010",
    580  => "1010101010101010",
    581  => "1010101010101010",
    582  => "1010101010101010",
    583  => "1010101010101010",
    584  => "1010101010101010",
    585  => "1010101010101010",
    586  => "1010101010101010",
    587  => "1010101010101010",
    588  => "1010101010101010",
    589  => "1010101010101010",
    590  => "1010101010101010",
    591  => "1010101010101010",
    592  => "1010101010101010",
    593  => "1010101010101010",
    594  => "1010101010101010",
    595  => "1010101010101010",
    596  => "1010101010101010",
    597  => "1010101010101010",
    598  => "1010101010101010",
    599  => "1010101010101010",
    600  => "1010101010101010",
    601  => "1010101010101010",
    602  => "1010101010101010",
    603  => "1010101010101010",
    604  => "1010101010101010",
    605  => "1010101010101010",
    606  => "1010101010101010",
    607  => "1010101010101010",
    608  => "1010101010101010",
    609  => "1010101010101010",
    610  => "1010101010101010",
    611  => "1010101010101010",
    612  => "1010101010101010",
    613  => "1010101010101010",
    614  => "1010101010101010",
    615  => "1010101010101010",
    616  => "1010101010101010",
    617  => "1010101010101010",
    618  => "1010101010101010",
    619  => "1010101010101010",
    620  => "1010101010101010",
    621  => "1010101010101010",
    622  => "1010101010101010",
    623  => "1010101010101010",
    624  => "1010101010101010",
    625  => "1010101010101010",
    626  => "1010101010101010",
    627  => "1010101010101010",
    628  => "1010101010101010",
    629  => "1010101010101010",
    630  => "1010101010101010",
    631  => "1010101010101010",
    632  => "1010101010101010",
    633  => "1010101010101010",
    634  => "1010101010101010",
    635  => "1010101010101010",
    636  => "1010101010101010",
    637  => "1010101010101010",
    638  => "1010101010101010",
    639  => "1010101010101010",
    640  => "1010101010101010",
    641  => "1010101010101010",
    642  => "1010101010101010",
    643  => "1010101010101010",
    644  => "1010101010101010",
    645  => "1010101010101010",
    646  => "1010101010101010",
    647  => "1010101010101010",
    648  => "1010101010101010",
    649  => "1010101010101010",
    650  => "1010101010101010",
    651  => "1010101010101010",
    652  => "1010101010101010",
    653  => "1010101010101010",
    654  => "1010101010101010",
    655  => "1010101010101010",
    656  => "1010101010101010",
    657  => "1010101010101010",
    658  => "1010101010101010",
    659  => "1010101010101010",
    660  => "1010101010101010",
    661  => "1010101010101010",
    662  => "1010101010101010",
    663  => "1010101010101010",
    664  => "1010101010101010",
    665  => "1010101010101010",
    666  => "1010101010101010",
    667  => "1010101010101010",
    668  => "1010101010101010",
    669  => "1010101010101010",
    670  => "1010101010101010",
    671  => "1010101010101010",
    672  => "1010101010101010",
    673  => "1010101010101010",
    674  => "1010101010101010",
    675  => "1010101010101010",
    676  => "1010101010101010",
    677  => "1010101010101010",
    678  => "1010101010101010",
    679  => "1010101010101010",
    680  => "1010101010101010",
    681  => "1010101010101010",
    682  => "1010101010101010",
    683  => "1010101010101010",
    684  => "1010101010101010",
    685  => "1010101010101010",
    686  => "1010101010101010",
    687  => "1010101010101010",
    688  => "1010101010101010",
    689  => "1010101010101010",
    690  => "1010101010101010",
    691  => "1010101010101010",
    692  => "1010101010101010",
    693  => "1010101010101010",
    694  => "1010101010101010",
    695  => "1010101010101010",
    696  => "1010101010101010",
    697  => "1010101010101010",
    698  => "1010101010101010",
    699  => "1010101010101010",
    700  => "1010101010101010",
    701  => "1010101010101010",
    702  => "1010101010101010",
    703  => "1010101010101010",
    704  => "1010101010101010",
    705  => "1010101010101010",
    706  => "1010101010101010",
    707  => "1010101010101010",
    708  => "1010101010101010",
    709  => "1010101010101010",
    710  => "1010101010101010",
    711  => "1010101010101010",
    712  => "1010101010101010",
    713  => "1010101010101010",
    714  => "1010101010101010",
    715  => "1010101010101010",
    716  => "1010101010101010",
    717  => "1010101010101010",
    718  => "1010101010101010",
    719  => "1010101010101010",
    720  => "1010101010101010",
    721  => "1010101010101010",
    722  => "1010101010101010",
    723  => "1010101010101010",
    724  => "1010101010101010",
    725  => "1010101010101010",
    726  => "1010101010101010",
    727  => "1010101010101010",
    728  => "1010101010101010",
    729  => "1010101010101010",
    730  => "1010101010101010",
    731  => "1010101010101010",
    732  => "1010101010101010",
    733  => "1010101010101010",
    734  => "1010101010101010",
    735  => "1010101010101010",
    736  => "1010101010101010",
    737  => "1010101010101010",
    738  => "1010101010101010",
    739  => "1010101010101010",
    740  => "1010101010101010",
    741  => "1010101010101010",
    742  => "1010101010101010",
    743  => "1010101010101010",
    744  => "1010101010101010",
    745  => "1010101010101010",
    746  => "1010101010101010",
    747  => "1010101010101010",
    748  => "1010101010101010",
    749  => "1010101010101010",
    750  => "1010101010101010",
    751  => "1010101010101010",
    752  => "1010101010101010",
    753  => "1010101010101010",
    754  => "1010101010101010",
    755  => "1010101010101010",
    756  => "1010101010101010",
    757  => "1010101010101010",
    758  => "1010101010101010",
    759  => "1010101010101010",
    760  => "1010101010101010",
    761  => "1010101010101010",
    762  => "1010101010101010",
    763  => "1010101010101010",
    764  => "1010101010101010",
    765  => "1010101010101010",
    766  => "1010101010101010",
    767  => "1010101010101010",
    768  => "1010101010101010",
    769  => "1010101010101010",
    770  => "1010101010101010",
    771  => "1010101010101010",
    772  => "1010101010101010",
    773  => "1010101010101010",
    774  => "1010101010101010",
    775  => "1010101010101010",
    776  => "1010101010101010",
    777  => "1010101010101010",
    778  => "1010101010101010",
    779  => "1010101010101010",
    780  => "1010101010101010",
    781  => "1010101010101010",
    782  => "1010101010101010",
    783  => "1010101010101010",
    784  => "1010101010101010",
    785  => "1010101010101010",
    786  => "1010101010101010",
    787  => "1010101010101010",
    788  => "1010101010101010",
    789  => "1010101010101010",
    790  => "1010101010101010",
    791  => "1010101010101010",
    792  => "1010101010101010",
    793  => "1010101010101010",
    794  => "1010101010101010",
    795  => "1010101010101010",
    796  => "1010101010101010",
    797  => "1010101010101010",
    798  => "1010101010101010",
    799  => "1010101010101010",
    800  => "1010101010101010",
    801  => "1010101010101010",
    802  => "1010101010101010",
    803  => "1010101010101010",
    804  => "1010101010101010",
    805  => "1010101010101010",
    806  => "1010101010101010",
    807  => "1010101010101010",
    808  => "1010101010101010",
    809  => "1010101010101010",
    810  => "1010101010101010",
    811  => "1010101010101010",
    812  => "1010101010101010",
    813  => "1010101010101010",
    814  => "1010101010101010",
    815  => "1010101010101010",
    816  => "1010101010101010",
    817  => "1010101010101010",
    818  => "1010101010101010",
    819  => "1010101010101010",
    820  => "1010101010101010",
    821  => "1010101010101010",
    822  => "1010101010101010",
    823  => "1010101010101010",
    824  => "1010101010101010",
    825  => "1010101010101010",
    826  => "1010101010101010",
    827  => "1010101010101010",
    828  => "1010101010101010",
    829  => "1010101010101010",
    830  => "1010101010101010",
    831  => "1010101010101010",
    832  => "1010101010101010",
    833  => "1010101010101010",
    834  => "1010101010101010",
    835  => "1010101010101010",
    836  => "1010101010101010",
    837  => "1010101010101010",
    838  => "1010101010101010",
    839  => "1010101010101010",
    840  => "1010101010101010",
    841  => "1010101010101010",
    842  => "1010101010101010",
    843  => "1010101010101010",
    844  => "1010101010101010",
    845  => "1010101010101010",
    846  => "1010101010101010",
    847  => "1010101010101010",
    848  => "1010101010101010",
    849  => "1010101010101010",
    850  => "1010101010101010",
    851  => "1010101010101010",
    852  => "1010101010101010",
    853  => "1010101010101010",
    854  => "1010101010101010",
    855  => "1010101010101010",
    856  => "1010101010101010",
    857  => "1010101010101010",
    858  => "1010101010101010",
    859  => "1010101010101010",
    860  => "1010101010101010",
    861  => "1010101010101010",
    862  => "1010101010101010",
    863  => "1010101010101010",
    864  => "1010101010101010",
    865  => "1010101010101010",
    866  => "1010101010101010",
    867  => "1010101010101010",
    868  => "1010101010101010",
    869  => "1010101010101010",
    870  => "1010101010101010",
    871  => "1010101010101010",
    872  => "1010101010101010",
    873  => "1010101010101010",
    874  => "1010101010101010",
    875  => "1010101010101010",
    876  => "1010101010101010",
    877  => "1010101010101010",
    878  => "1010101010101010",
    879  => "1010101010101010",
    880  => "1010101010101010",
    881  => "1010101010101010",
    882  => "1010101010101010",
    883  => "1010101010101010",
    884  => "1010101010101010",
    885  => "1010101010101010",
    886  => "1010101010101010",
    887  => "1010101010101010",
    888  => "1010101010101010",
    889  => "1010101010101010",
    890  => "1010101010101010",
    891  => "1010101010101010",
    892  => "1010101010101010",
    893  => "1010101010101010",
    894  => "1010101010101010",
    895  => "1010101010101010",
    896  => "1010101010101010",
    897  => "1010101010101010",
    898  => "1010101010101010",
    899  => "1010101010101010",
    900  => "1010101010101010",
    901  => "1010101010101010",
    902  => "1010101010101010",
    903  => "1010101010101010",
    904  => "1010101010101010",
    905  => "1010101010101010",
    906  => "1010101010101010",
    907  => "1010101010101010",
    908  => "1010101010101010",
    909  => "1010101010101010",
    910  => "1010101010101010",
    911  => "1010101010101010",
    912  => "1010101010101010",
    913  => "1010101010101010",
    914  => "1010101010101010",
    915  => "1010101010101010",
    916  => "1010101010101010",
    917  => "1010101010101010",
    918  => "1010101010101010",
    919  => "1010101010101010",
    920  => "1010101010101010",
    921  => "1010101010101010",
    922  => "1010101010101010",
    923  => "1010101010101010",
    924  => "1010101010101010",
    925  => "1010101010101010",
    926  => "1010101010101010",
    927  => "1010101010101010",
    928  => "1010101010101010",
    929  => "1010101010101010",
    930  => "1010101010101010",
    931  => "1010101010101010",
    932  => "1010101010101010",
    933  => "1010101010101010",
    934  => "1010101010101010",
    935  => "1010101010101010",
    936  => "1010101010101010",
    937  => "1010101010101010",
    938  => "1010101010101010",
    939  => "1010101010101010",
    940  => "1010101010101010",
    941  => "1010101010101010",
    942  => "1010101010101010",
    943  => "1010101010101010",
    944  => "1010101010101010",
    945  => "1010101010101010",
    946  => "1010101010101010",
    947  => "1010101010101010",
    948  => "1010101010101010",
    949  => "1010101010101010",
    950  => "1010101010101010",
    951  => "1010101010101010",
    952  => "1010101010101010",
    953  => "1010101010101010",
    954  => "1010101010101010",
    955  => "1010101010101010",
    956  => "1010101010101010",
    957  => "1010101010101010",
    958  => "1010101010101010",
    959  => "1010101010101010",
    960  => "1010101010101010",
    961  => "1010101010101010",
    962  => "1010101010101010",
    963  => "1010101010101010",
    964  => "1010101010101010",
    965  => "1010101010101010",
    966  => "1010101010101010",
    967  => "1010101010101010",
    968  => "1010101010101010",
    969  => "1010101010101010",
    970  => "1010101010101010",
    971  => "1010101010101010",
    972  => "1010101010101010",
    973  => "1010101010101010",
    974  => "1010101010101010",
    975  => "1010101010101010",
    976  => "1010101010101010",
    977  => "1010101010101010",
    978  => "1010101010101010",
    979  => "1010101010101010",
    980  => "1010101010101010",
    981  => "1010101010101010",
    982  => "1010101010101010",
    983  => "1010101010101010",
    984  => "1010101010101010",
    985  => "1010101010101010",
    986  => "1010101010101010",
    987  => "1010101010101010",
    988  => "1010101010101010",
    989  => "1010101010101010",
    990  => "1010101010101010",
    991  => "1010101010101010",
    992  => "1010101010101010",
    993  => "1010101010101010",
    994  => "1010101010101010",
    995  => "1010101010101010",
    996  => "1010101010101010",
    997  => "1010101010101010",
    998  => "1010101010101010",
    999  => "1010101010101010",
    1000 => "1010101010101010",
    1001 => "1010101010101010",
    1002 => "1010101010101010",
    1003 => "1010101010101010",
    1004 => "1010101010101010",
    1005 => "1010101010101010",
    1006 => "1010101010101010",
    1007 => "1010101010101010",
    1008 => "1010101010101010",
    1009 => "1010101010101010",
    1010 => "1010101010101010",
    1011 => "1010101010101010",
    1012 => "1010101010101010",
    1013 => "1010101010101010",
    1014 => "1010101010101010",
    1015 => "1010101010101010",
    1016 => "1010101010101010",
    1017 => "1010101010101010",
    1018 => "1010101010101010",
    1019 => "1010101010101010",
    1020 => "1010101010101010",
    1021 => "1010101010101010",
    1022 => "1010101010101010",
    1023 => "1010101010101010"
    );

end mem_buffer;