library ieee;
use ieee.std_logic_1164.all;

package svnr_memory_image is
  constant address_size : integer := 10;  -- ram_adddress breite
  type mem_type is array (0 to (2**address_size)-1) of std_logic_vector(15 downto 0);

  constant mem_init_image : mem_type := (
      0 => x"4820",
      1 => x"0000",
      2 => x"0000",
      3 => x"0000",
      4 => x"0000",
      5 => x"0000",
      6 => x"5555",
      7 => x"0000",
      8 => x"0000",
      9 => x"0000",
     10 => x"0000",
     11 => x"0000",
     12 => x"0000",
     13 => x"0000",
     14 => x"0000",
     15 => x"0000",
     16 => x"0000",
     17 => x"0003",
     18 => x"000f",
     19 => x"0005",
     20 => x"0000",
     21 => x"0000",
     22 => x"0000",
     23 => x"0000",
     24 => x"0000",
     25 => x"0000",
     26 => x"0000",
     27 => x"0000",
     28 => x"0000",
     29 => x"0000",
     30 => x"0000",
     31 => x"0000",
     32 => x"1112",
     33 => x"3111",
     34 => x"582a",
     35 => x"1113",
     36 => x"3900",
     37 => x"2813",
     38 => x"482f",
     39 => x"0000",
     40 => x"0000",
     41 => x"0000",
     42 => x"1113",
     43 => x"3800",
     44 => x"2813",
     45 => x"1000",
     46 => x"1000",
     47 => x"482f",
     48 => x"0000",
     49 => x"0000",
     50 => x"0000",
     51 => x"0000",
     52 => x"0000",
     53 => x"0000",
     54 => x"0000",
     55 => x"0000",
     56 => x"0000",
     57 => x"0000",
     58 => x"0000",
     59 => x"0000",
     60 => x"0000",
     61 => x"0000",
     62 => x"0000",
     63 => x"0000",
     64 => x"0000",
     65 => x"0000",
     66 => x"0000",
     67 => x"0000",
     68 => x"0000",
     69 => x"0000",
     70 => x"0000",
     71 => x"0000",
     72 => x"0000",
     73 => x"0000",
     74 => x"0000",
     75 => x"0000",
     76 => x"0000",
     77 => x"0000",
     78 => x"0000",
     79 => x"0000",
     80 => x"0000",
     81 => x"0000",
     82 => x"0000",
     83 => x"0000",
     84 => x"0000",
     85 => x"0000",
     86 => x"0000",
     87 => x"0000",
     88 => x"0000",
     89 => x"0000",
     90 => x"0000",
     91 => x"0000",
     92 => x"0000",
     93 => x"0000",
     94 => x"0000",
     95 => x"0000",
     96 => x"0000",
     97 => x"0000",
     98 => x"0000",
     99 => x"0000",
    100 => x"0000",
    101 => x"0000",
    102 => x"0000",
    103 => x"0000",
    104 => x"0000",
    105 => x"0000",
    106 => x"0000",
    107 => x"0000",
    108 => x"0000",
    109 => x"0000",
    110 => x"0000",
    111 => x"0000",
    112 => x"0000",
    113 => x"0000",
    114 => x"0000",
    115 => x"0000",
    116 => x"0000",
    117 => x"0000",
    118 => x"0000",
    119 => x"0000",
    120 => x"0000",
    121 => x"0000",
    122 => x"0000",
    123 => x"0000",
    124 => x"0000",
    125 => x"0000",
    126 => x"0000",
    127 => x"0000",
    128 => x"0000",
    129 => x"0000",
    130 => x"0000",
    131 => x"0000",
    132 => x"0000",
    133 => x"0000",
    134 => x"0000",
    135 => x"0000",
    136 => x"0000",
    137 => x"0000",
    138 => x"0000",
    139 => x"0000",
    140 => x"0000",
    141 => x"0000",
    142 => x"0000",
    143 => x"0000",
    144 => x"0000",
    145 => x"0000",
    146 => x"0000",
    147 => x"0000",
    148 => x"0000",
    149 => x"0000",
    150 => x"0000",
    151 => x"0000",
    152 => x"0000",
    153 => x"0000",
    154 => x"0000",
    155 => x"0000",
    156 => x"0000",
    157 => x"0000",
    158 => x"0000",
    159 => x"0000",
    160 => x"0000",
    161 => x"0000",
    162 => x"0000",
    163 => x"0000",
    164 => x"0000",
    165 => x"0000",
    166 => x"0000",
    167 => x"0000",
    168 => x"0000",
    169 => x"0000",
    170 => x"0000",
    171 => x"0000",
    172 => x"0000",
    173 => x"0000",
    174 => x"0000",
    175 => x"0000",
    176 => x"0000",
    177 => x"0000",
    178 => x"0000",
    179 => x"0000",
    180 => x"0000",
    181 => x"0000",
    182 => x"0000",
    183 => x"0000",
    184 => x"0000",
    185 => x"0000",
    186 => x"0000",
    187 => x"0000",
    188 => x"0000",
    189 => x"0000",
    190 => x"0000",
    191 => x"0000",
    192 => x"0000",
    193 => x"0000",
    194 => x"0000",
    195 => x"0000",
    196 => x"0000",
    197 => x"0000",
    198 => x"0000",
    199 => x"0000",
    200 => x"0000",
    201 => x"0000",
    202 => x"0000",
    203 => x"0000",
    204 => x"0000",
    205 => x"0000",
    206 => x"0000",
    207 => x"0000",
    208 => x"0000",
    209 => x"0000",
    210 => x"0000",
    211 => x"0000",
    212 => x"0000",
    213 => x"0000",
    214 => x"0000",
    215 => x"0000",
    216 => x"0000",
    217 => x"0000",
    218 => x"0000",
    219 => x"0000",
    220 => x"0000",
    221 => x"0000",
    222 => x"0000",
    223 => x"0000",
    224 => x"0000",
    225 => x"0000",
    226 => x"0000",
    227 => x"0000",
    228 => x"0000",
    229 => x"0000",
    230 => x"0000",
    231 => x"0000",
    232 => x"0000",
    233 => x"0000",
    234 => x"0000",
    235 => x"0000",
    236 => x"0000",
    237 => x"0000",
    238 => x"0000",
    239 => x"0000",
    240 => x"0000",
    241 => x"0000",
    242 => x"0000",
    243 => x"0000",
    244 => x"0000",
    245 => x"0000",
    246 => x"0000",
    247 => x"0000",
    248 => x"0000",
    249 => x"0000",
    250 => x"0000",
    251 => x"0000",
    252 => x"0000",
    253 => x"0000",
    254 => x"0000",
    255 => x"0000",
    256 => x"0000",
    257 => x"0000",
    258 => x"0000",
    259 => x"0000",
    260 => x"0000",
    261 => x"0000",
    262 => x"0000",
    263 => x"0000",
    264 => x"0000",
    265 => x"0000",
    266 => x"0000",
    267 => x"0000",
    268 => x"0000",
    269 => x"0000",
    270 => x"0000",
    271 => x"0000",
    272 => x"0000",
    273 => x"0000",
    274 => x"0000",
    275 => x"0000",
    276 => x"0000",
    277 => x"0000",
    278 => x"0000",
    279 => x"0000",
    280 => x"0000",
    281 => x"0000",
    282 => x"0000",
    283 => x"0000",
    284 => x"0000",
    285 => x"0000",
    286 => x"0000",
    287 => x"0000",
    288 => x"0000",
    289 => x"0000",
    290 => x"0000",
    291 => x"0000",
    292 => x"0000",
    293 => x"0000",
    294 => x"0000",
    295 => x"0000",
    296 => x"0000",
    297 => x"0000",
    298 => x"0000",
    299 => x"0000",
    300 => x"0000",
    301 => x"0000",
    302 => x"0000",
    303 => x"0000",
    304 => x"0000",
    305 => x"0000",
    306 => x"0000",
    307 => x"0000",
    308 => x"0000",
    309 => x"0000",
    310 => x"0000",
    311 => x"0000",
    312 => x"0000",
    313 => x"0000",
    314 => x"0000",
    315 => x"0000",
    316 => x"0000",
    317 => x"0000",
    318 => x"0000",
    319 => x"0000",
    320 => x"0000",
    321 => x"0000",
    322 => x"0000",
    323 => x"0000",
    324 => x"0000",
    325 => x"0000",
    326 => x"0000",
    327 => x"0000",
    328 => x"0000",
    329 => x"0000",
    330 => x"0000",
    331 => x"0000",
    332 => x"0000",
    333 => x"0000",
    334 => x"0000",
    335 => x"0000",
    336 => x"0000",
    337 => x"0000",
    338 => x"0000",
    339 => x"0000",
    340 => x"0000",
    341 => x"0000",
    342 => x"0000",
    343 => x"0000",
    344 => x"0000",
    345 => x"0000",
    346 => x"0000",
    347 => x"0000",
    348 => x"0000",
    349 => x"0000",
    350 => x"0000",
    351 => x"0000",
    352 => x"0000",
    353 => x"0000",
    354 => x"0000",
    355 => x"0000",
    356 => x"0000",
    357 => x"0000",
    358 => x"0000",
    359 => x"0000",
    360 => x"0000",
    361 => x"0000",
    362 => x"0000",
    363 => x"0000",
    364 => x"0000",
    365 => x"0000",
    366 => x"0000",
    367 => x"0000",
    368 => x"0000",
    369 => x"0000",
    370 => x"0000",
    371 => x"0000",
    372 => x"0000",
    373 => x"0000",
    374 => x"0000",
    375 => x"0000",
    376 => x"0000",
    377 => x"0000",
    378 => x"0000",
    379 => x"0000",
    380 => x"0000",
    381 => x"0000",
    382 => x"0000",
    383 => x"0000",
    384 => x"0000",
    385 => x"0000",
    386 => x"0000",
    387 => x"0000",
    388 => x"0000",
    389 => x"0000",
    390 => x"0000",
    391 => x"0000",
    392 => x"0000",
    393 => x"0000",
    394 => x"0000",
    395 => x"0000",
    396 => x"0000",
    397 => x"0000",
    398 => x"0000",
    399 => x"0000",
    400 => x"0000",
    401 => x"0000",
    402 => x"0000",
    403 => x"0000",
    404 => x"0000",
    405 => x"0000",
    406 => x"0000",
    407 => x"0000",
    408 => x"0000",
    409 => x"0000",
    410 => x"0000",
    411 => x"0000",
    412 => x"0000",
    413 => x"0000",
    414 => x"0000",
    415 => x"0000",
    416 => x"0000",
    417 => x"0000",
    418 => x"0000",
    419 => x"0000",
    420 => x"0000",
    421 => x"0000",
    422 => x"0000",
    423 => x"0000",
    424 => x"0000",
    425 => x"0000",
    426 => x"0000",
    427 => x"0000",
    428 => x"0000",
    429 => x"0000",
    430 => x"0000",
    431 => x"0000",
    432 => x"0000",
    433 => x"0000",
    434 => x"0000",
    435 => x"0000",
    436 => x"0000",
    437 => x"0000",
    438 => x"0000",
    439 => x"0000",
    440 => x"0000",
    441 => x"0000",
    442 => x"0000",
    443 => x"0000",
    444 => x"0000",
    445 => x"0000",
    446 => x"0000",
    447 => x"0000",
    448 => x"0000",
    449 => x"0000",
    450 => x"0000",
    451 => x"0000",
    452 => x"0000",
    453 => x"0000",
    454 => x"0000",
    455 => x"0000",
    456 => x"0000",
    457 => x"0000",
    458 => x"0000",
    459 => x"0000",
    460 => x"0000",
    461 => x"0000",
    462 => x"0000",
    463 => x"0000",
    464 => x"0000",
    465 => x"0000",
    466 => x"0000",
    467 => x"0000",
    468 => x"0000",
    469 => x"0000",
    470 => x"0000",
    471 => x"0000",
    472 => x"0000",
    473 => x"0000",
    474 => x"0000",
    475 => x"0000",
    476 => x"0000",
    477 => x"0000",
    478 => x"0000",
    479 => x"0000",
    480 => x"0000",
    481 => x"0000",
    482 => x"0000",
    483 => x"0000",
    484 => x"0000",
    485 => x"0000",
    486 => x"0000",
    487 => x"0000",
    488 => x"0000",
    489 => x"0000",
    490 => x"0000",
    491 => x"0000",
    492 => x"0000",
    493 => x"0000",
    494 => x"0000",
    495 => x"0000",
    496 => x"0000",
    497 => x"0000",
    498 => x"0000",
    499 => x"0000",
    500 => x"0000",
    501 => x"0000",
    502 => x"0000",
    503 => x"0000",
    504 => x"0000",
    505 => x"0000",
    506 => x"0000",
    507 => x"0000",
    508 => x"0000",
    509 => x"0000",
    510 => x"0000",
    511 => x"0000",
    512 => x"0000",
    513 => x"0000",
    514 => x"0000",
    515 => x"0000",
    516 => x"0000",
    517 => x"0000",
    518 => x"0000",
    519 => x"0000",
    520 => x"0000",
    521 => x"0000",
    522 => x"0000",
    523 => x"0000",
    524 => x"0000",
    525 => x"0000",
    526 => x"0000",
    527 => x"0000",
    528 => x"0000",
    529 => x"0000",
    530 => x"0000",
    531 => x"0000",
    532 => x"0000",
    533 => x"0000",
    534 => x"0000",
    535 => x"0000",
    536 => x"0000",
    537 => x"0000",
    538 => x"0000",
    539 => x"0000",
    540 => x"0000",
    541 => x"0000",
    542 => x"0000",
    543 => x"0000",
    544 => x"0000",
    545 => x"0000",
    546 => x"0000",
    547 => x"0000",
    548 => x"0000",
    549 => x"0000",
    550 => x"0000",
    551 => x"0000",
    552 => x"0000",
    553 => x"0000",
    554 => x"0000",
    555 => x"0000",
    556 => x"0000",
    557 => x"0000",
    558 => x"0000",
    559 => x"0000",
    560 => x"0000",
    561 => x"0000",
    562 => x"0000",
    563 => x"0000",
    564 => x"0000",
    565 => x"0000",
    566 => x"0000",
    567 => x"0000",
    568 => x"0000",
    569 => x"0000",
    570 => x"0000",
    571 => x"0000",
    572 => x"0000",
    573 => x"0000",
    574 => x"0000",
    575 => x"0000",
    576 => x"0000",
    577 => x"0000",
    578 => x"0000",
    579 => x"0000",
    580 => x"0000",
    581 => x"0000",
    582 => x"0000",
    583 => x"0000",
    584 => x"0000",
    585 => x"0000",
    586 => x"0000",
    587 => x"0000",
    588 => x"0000",
    589 => x"0000",
    590 => x"0000",
    591 => x"0000",
    592 => x"0000",
    593 => x"0000",
    594 => x"0000",
    595 => x"0000",
    596 => x"0000",
    597 => x"0000",
    598 => x"0000",
    599 => x"0000",
    600 => x"0000",
    601 => x"0000",
    602 => x"0000",
    603 => x"0000",
    604 => x"0000",
    605 => x"0000",
    606 => x"0000",
    607 => x"0000",
    608 => x"0000",
    609 => x"0000",
    610 => x"0000",
    611 => x"0000",
    612 => x"0000",
    613 => x"0000",
    614 => x"0000",
    615 => x"0000",
    616 => x"0000",
    617 => x"0000",
    618 => x"0000",
    619 => x"0000",
    620 => x"0000",
    621 => x"0000",
    622 => x"0000",
    623 => x"0000",
    624 => x"0000",
    625 => x"0000",
    626 => x"0000",
    627 => x"0000",
    628 => x"0000",
    629 => x"0000",
    630 => x"0000",
    631 => x"0000",
    632 => x"0000",
    633 => x"0000",
    634 => x"0000",
    635 => x"0000",
    636 => x"0000",
    637 => x"0000",
    638 => x"0000",
    639 => x"0000",
    640 => x"0000",
    641 => x"0000",
    642 => x"0000",
    643 => x"0000",
    644 => x"0000",
    645 => x"0000",
    646 => x"0000",
    647 => x"0000",
    648 => x"0000",
    649 => x"0000",
    650 => x"0000",
    651 => x"0000",
    652 => x"0000",
    653 => x"0000",
    654 => x"0000",
    655 => x"0000",
    656 => x"0000",
    657 => x"0000",
    658 => x"0000",
    659 => x"0000",
    660 => x"0000",
    661 => x"0000",
    662 => x"0000",
    663 => x"0000",
    664 => x"0000",
    665 => x"0000",
    666 => x"0000",
    667 => x"0000",
    668 => x"0000",
    669 => x"0000",
    670 => x"0000",
    671 => x"0000",
    672 => x"0000",
    673 => x"0000",
    674 => x"0000",
    675 => x"0000",
    676 => x"0000",
    677 => x"0000",
    678 => x"0000",
    679 => x"0000",
    680 => x"0000",
    681 => x"0000",
    682 => x"0000",
    683 => x"0000",
    684 => x"0000",
    685 => x"0000",
    686 => x"0000",
    687 => x"0000",
    688 => x"0000",
    689 => x"0000",
    690 => x"0000",
    691 => x"0000",
    692 => x"0000",
    693 => x"0000",
    694 => x"0000",
    695 => x"0000",
    696 => x"0000",
    697 => x"0000",
    698 => x"0000",
    699 => x"0000",
    700 => x"0000",
    701 => x"0000",
    702 => x"0000",
    703 => x"0000",
    704 => x"0000",
    705 => x"0000",
    706 => x"0000",
    707 => x"0000",
    708 => x"0000",
    709 => x"0000",
    710 => x"0000",
    711 => x"0000",
    712 => x"0000",
    713 => x"0000",
    714 => x"0000",
    715 => x"0000",
    716 => x"0000",
    717 => x"0000",
    718 => x"0000",
    719 => x"0000",
    720 => x"0000",
    721 => x"0000",
    722 => x"0000",
    723 => x"0000",
    724 => x"0000",
    725 => x"0000",
    726 => x"0000",
    727 => x"0000",
    728 => x"0000",
    729 => x"0000",
    730 => x"0000",
    731 => x"0000",
    732 => x"0000",
    733 => x"0000",
    734 => x"0000",
    735 => x"0000",
    736 => x"0000",
    737 => x"0000",
    738 => x"0000",
    739 => x"0000",
    740 => x"0000",
    741 => x"0000",
    742 => x"0000",
    743 => x"0000",
    744 => x"0000",
    745 => x"0000",
    746 => x"0000",
    747 => x"0000",
    748 => x"0000",
    749 => x"0000",
    750 => x"0000",
    751 => x"0000",
    752 => x"0000",
    753 => x"0000",
    754 => x"0000",
    755 => x"0000",
    756 => x"0000",
    757 => x"0000",
    758 => x"0000",
    759 => x"0000",
    760 => x"0000",
    761 => x"0000",
    762 => x"0000",
    763 => x"0000",
    764 => x"0000",
    765 => x"0000",
    766 => x"0000",
    767 => x"0000",
    768 => x"0000",
    769 => x"0000",
    770 => x"0000",
    771 => x"0000",
    772 => x"0000",
    773 => x"0000",
    774 => x"0000",
    775 => x"0000",
    776 => x"0000",
    777 => x"0000",
    778 => x"0000",
    779 => x"0000",
    780 => x"0000",
    781 => x"0000",
    782 => x"0000",
    783 => x"0000",
    784 => x"0000",
    785 => x"0000",
    786 => x"0000",
    787 => x"0000",
    788 => x"0000",
    789 => x"0000",
    790 => x"0000",
    791 => x"0000",
    792 => x"0000",
    793 => x"0000",
    794 => x"0000",
    795 => x"0000",
    796 => x"0000",
    797 => x"0000",
    798 => x"0000",
    799 => x"0000",
    800 => x"0000",
    801 => x"0000",
    802 => x"0000",
    803 => x"0000",
    804 => x"0000",
    805 => x"0000",
    806 => x"0000",
    807 => x"0000",
    808 => x"0000",
    809 => x"0000",
    810 => x"0000",
    811 => x"0000",
    812 => x"0000",
    813 => x"0000",
    814 => x"0000",
    815 => x"0000",
    816 => x"0000",
    817 => x"0000",
    818 => x"0000",
    819 => x"0000",
    820 => x"0000",
    821 => x"0000",
    822 => x"0000",
    823 => x"0000",
    824 => x"0000",
    825 => x"0000",
    826 => x"0000",
    827 => x"0000",
    828 => x"0000",
    829 => x"0000",
    830 => x"0000",
    831 => x"0000",
    832 => x"0000",
    833 => x"0000",
    834 => x"0000",
    835 => x"0000",
    836 => x"0000",
    837 => x"0000",
    838 => x"0000",
    839 => x"0000",
    840 => x"0000",
    841 => x"0000",
    842 => x"0000",
    843 => x"0000",
    844 => x"0000",
    845 => x"0000",
    846 => x"0000",
    847 => x"0000",
    848 => x"0000",
    849 => x"0000",
    850 => x"0000",
    851 => x"0000",
    852 => x"0000",
    853 => x"0000",
    854 => x"0000",
    855 => x"0000",
    856 => x"0000",
    857 => x"0000",
    858 => x"0000",
    859 => x"0000",
    860 => x"0000",
    861 => x"0000",
    862 => x"0000",
    863 => x"0000",
    864 => x"0000",
    865 => x"0000",
    866 => x"0000",
    867 => x"0000",
    868 => x"0000",
    869 => x"0000",
    870 => x"0000",
    871 => x"0000",
    872 => x"0000",
    873 => x"0000",
    874 => x"0000",
    875 => x"0000",
    876 => x"0000",
    877 => x"0000",
    878 => x"0000",
    879 => x"0000",
    880 => x"0000",
    881 => x"0000",
    882 => x"0000",
    883 => x"0000",
    884 => x"0000",
    885 => x"0000",
    886 => x"0000",
    887 => x"0000",
    888 => x"0000",
    889 => x"0000",
    890 => x"0000",
    891 => x"0000",
    892 => x"0000",
    893 => x"0000",
    894 => x"0000",
    895 => x"0000",
    896 => x"0000",
    897 => x"0000",
    898 => x"0000",
    899 => x"0000",
    900 => x"0000",
    901 => x"0000",
    902 => x"0000",
    903 => x"0000",
    904 => x"0000",
    905 => x"0000",
    906 => x"0000",
    907 => x"0000",
    908 => x"0000",
    909 => x"0000",
    910 => x"0000",
    911 => x"0000",
    912 => x"0000",
    913 => x"0000",
    914 => x"0000",
    915 => x"0000",
    916 => x"0000",
    917 => x"0000",
    918 => x"0000",
    919 => x"0000",
    920 => x"0000",
    921 => x"0000",
    922 => x"0000",
    923 => x"0000",
    924 => x"0000",
    925 => x"0000",
    926 => x"0000",
    927 => x"0000",
    928 => x"0000",
    929 => x"0000",
    930 => x"0000",
    931 => x"0000",
    932 => x"0000",
    933 => x"0000",
    934 => x"0000",
    935 => x"0000",
    936 => x"0000",
    937 => x"0000",
    938 => x"0000",
    939 => x"0000",
    940 => x"0000",
    941 => x"0000",
    942 => x"0000",
    943 => x"0000",
    944 => x"0000",
    945 => x"0000",
    946 => x"0000",
    947 => x"0000",
    948 => x"0000",
    949 => x"0000",
    950 => x"0000",
    951 => x"0000",
    952 => x"0000",
    953 => x"0000",
    954 => x"0000",
    955 => x"0000",
    956 => x"0000",
    957 => x"0000",
    958 => x"0000",
    959 => x"0000",
    960 => x"0000",
    961 => x"0000",
    962 => x"0000",
    963 => x"0000",
    964 => x"0000",
    965 => x"0000",
    966 => x"0000",
    967 => x"0000",
    968 => x"0000",
    969 => x"0000",
    970 => x"0000",
    971 => x"0000",
    972 => x"0000",
    973 => x"0000",
    974 => x"0000",
    975 => x"0000",
    976 => x"0000",
    977 => x"0000",
    978 => x"0000",
    979 => x"0000",
    980 => x"0000",
    981 => x"0000",
    982 => x"0000",
    983 => x"0000",
    984 => x"0000",
    985 => x"0000",
    986 => x"0000",
    987 => x"0000",
    988 => x"0000",
    989 => x"0000",
    990 => x"0000",
    991 => x"0000",
    992 => x"0000",
    993 => x"0000",
    994 => x"0000",
    995 => x"0000",
    996 => x"0000",
    997 => x"0000",
    998 => x"0000",
    999 => x"0000",
    1000 => x"0000",
    1001 => x"0000",
    1002 => x"0000",
    1003 => x"0000",
    1004 => x"0000",
    1005 => x"0000",
    1006 => x"0000",
    1007 => x"0000",
    1008 => x"0000",
    1009 => x"0000",
    1010 => x"0000",
    1011 => x"0000",
    1012 => x"0000",
    1013 => x"0000",
    1014 => x"0000",
    1015 => x"0000",
    1016 => x"0000",
    1017 => x"0000",
    1018 => x"0000",
    1019 => x"0000",
    1020 => x"0000",
    1021 => x"0000",
    1022 => x"0000",
    1023 => x"0000"
    );

end svnr_memory_image;
